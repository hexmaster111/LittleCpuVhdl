module LittleCpu (
    i_clk,
    i_rst
);




    
endmodule;
