localparam //Cpu Opcodes 
    OP_add = 4'd0,
    OP_xor = 4'd1;

localparam //alu opcodes
    ALU_XOR = 1,
    ALU_ADD = 0;
